LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY cont5 IS
	PORT(clock,enable,reset : IN STD_LOGIC;
		 sal : OUT STD_LOGIC;
		 Q : Buffer STD_LOGIC_VECTOR (3 downto 0));
END cont5;

ARCHITECTURE sol OF cont5 IS
BEGIN

	PROCESS(clock,reset)
	BEGIN
		if reset='0' then Q<="0000";sal<='0';
  		elsif (clock'event and clock='1') then
			if enable='1' then
				if (Q="0101") then Q<="0000";sal<='1';
				else Q<=Q+1;sal<='0';
				end if;
			end if;
		end if;
	END PROCESS;
END sol;